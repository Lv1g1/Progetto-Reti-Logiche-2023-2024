-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb_max_dimensione is
end tb_max_dimensione;

architecture tb_max_dimensione_arch of tb_max_dimensione is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    constant SCENARIO_LENGTH : integer := 1023;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

    signal scenario_input : scenario_type := (176, 0, 66, 0, 159, 0, 63, 0, 164, 0, 33, 0, 114, 0, 93, 0, 199, 0, 84, 0, 160, 0, 237, 0, 44, 0, 21, 0, 80, 0, 0, 0, 115, 0, 113, 0, 229, 0, 132, 0, 171, 0, 6, 0, 202, 0, 44, 0, 173, 0, 144, 0, 212, 0, 51, 0, 15, 0, 173, 0, 140, 0, 126, 0, 12, 0, 252, 0, 195, 0, 254, 0, 249, 0, 215, 0, 17, 0, 180, 0, 33, 0, 163, 0, 186, 0, 207, 0, 16, 0, 200, 0, 157, 0, 48, 0, 214, 0, 87, 0, 118, 0, 71, 0, 18, 0, 13, 0, 13, 0, 177, 0, 80, 0, 56, 0, 20, 0, 73, 0, 24, 0, 29, 0, 214, 0, 82, 0, 191, 0, 0, 0, 195, 0, 254, 0, 40, 0, 222, 0, 170, 0, 123, 0, 215, 0, 189, 0, 146, 0, 132, 0, 71, 0, 208, 0, 203, 0, 193, 0, 234, 0, 1, 0, 245, 0, 117, 0, 23, 0, 0, 0, 113, 0, 121, 0, 26, 0, 79, 0, 223, 0, 137, 0, 209, 0, 64, 0, 252, 0, 9, 0, 13, 0, 226, 0, 2, 0, 42, 0, 174, 0, 122, 0, 219, 0, 219, 0, 33, 0, 239, 0, 179, 0, 122, 0, 64, 0, 13, 0, 72, 0, 125, 0, 205, 0, 162, 0, 59, 0, 113, 0, 43, 0, 63, 0, 224, 0, 14, 0, 94, 0, 33, 0, 66, 0, 20, 0, 49, 0, 160, 0, 52, 0, 34, 0, 9, 0, 253, 0, 27, 0, 14, 0, 135, 0, 109, 0, 204, 0, 121, 0, 237, 0, 171, 0, 173, 0, 112, 0, 133, 0, 247, 0, 81, 0, 35, 0, 73, 0, 129, 0, 152, 0, 193, 0, 92, 0, 74, 0, 45, 0, 12, 0, 54, 0, 36, 0, 224, 0, 93, 0, 84, 0, 37, 0, 39, 0, 188, 0, 245, 0, 112, 0, 239, 0, 243, 0, 14, 0, 135, 0, 225, 0, 78, 0, 103, 0, 34, 0, 0, 0, 6, 0, 81, 0, 254, 0, 11, 0, 121, 0, 217, 0, 119, 0, 39, 0, 130, 0, 190, 0, 18, 0, 145, 0, 190, 0, 72, 0, 251, 0, 222, 0, 172, 0, 200, 0, 136, 0, 120, 0, 37, 0, 86, 0, 125, 0, 160, 0, 94, 0, 222, 0, 146, 0, 146, 0, 221, 0, 66, 0, 247, 0, 129, 0, 150, 0, 188, 0, 67, 0, 19, 0, 128, 0, 158, 0, 146, 0, 206, 0, 99, 0, 48, 0, 220, 0, 3, 0, 173, 0, 67, 0, 3, 0, 126, 0, 203, 0, 234, 0, 81, 0, 0, 0, 11, 0, 227, 0, 162, 0, 38, 0, 156, 0, 17, 0, 95, 0, 202, 0, 209, 0, 145, 0, 134, 0, 57, 0, 136, 0, 159, 0, 103, 0, 37, 0, 12, 0, 209, 0, 187, 0, 219, 0, 177, 0, 244, 0, 121, 0, 220, 0, 59, 0, 91, 0, 155, 0, 119, 0, 58, 0, 115, 0, 235, 0, 67, 0, 79, 0, 28, 0, 107, 0, 7, 0, 120, 0, 7, 0, 131, 0, 204, 0, 77, 0, 158, 0, 201, 0, 120, 0, 168, 0, 110, 0, 81, 0, 238, 0, 189, 0, 188, 0, 67, 0, 51, 0, 185, 0, 153, 0, 219, 0, 35, 0, 192, 0, 149, 0, 110, 0, 97, 0, 227, 0, 67, 0, 245, 0, 138, 0, 99, 0, 7, 0, 189, 0, 51, 0, 185, 0, 0, 0, 235, 0, 56, 0, 245, 0, 46, 0, 233, 0, 54, 0, 179, 0, 95, 0, 221, 0, 78, 0, 253, 0, 183, 0, 229, 0, 119, 0, 67, 0, 172, 0, 58, 0, 16, 0, 166, 0, 150, 0, 192, 0, 54, 0, 234, 0, 176, 0, 96, 0, 175, 0, 106, 0, 181, 0, 48, 0, 85, 0, 202, 0, 154, 0, 151, 0, 66, 0, 104, 0, 28, 0, 244, 0, 76, 0, 183, 0, 254, 0, 150, 0, 117, 0, 243, 0, 153, 0, 65, 0, 184, 0, 30, 0, 177, 0, 245, 0, 225, 0, 255, 0, 173, 0, 127, 0, 163, 0, 204, 0, 59, 0, 68, 0, 76, 0, 181, 0, 96, 0, 131, 0, 14, 0, 242, 0, 35, 0, 31, 0, 195, 0, 145, 0, 153, 0, 12, 0, 180, 0, 175, 0, 248, 0, 73, 0, 100, 0, 4, 0, 186, 0, 14, 0, 170, 0, 194, 0, 102, 0, 118, 0, 252, 0, 191, 0, 175, 0, 245, 0, 182, 0, 75, 0, 210, 0, 41, 0, 177, 0, 101, 0, 149, 0, 9, 0, 119, 0, 30, 0, 49, 0, 119, 0, 164, 0, 118, 0, 245, 0, 105, 0, 92, 0, 201, 0, 175, 0, 167, 0, 224, 0, 99, 0, 14, 0, 63, 0, 104, 0, 189, 0, 174, 0, 84, 0, 160, 0, 206, 0, 4, 0, 20, 0, 173, 0, 187, 0, 82, 0, 46, 0, 234, 0, 217, 0, 20, 0, 47, 0, 8, 0, 119, 0, 31, 0, 198, 0, 25, 0, 170, 0, 139, 0, 218, 0, 4, 0, 207, 0, 65, 0, 222, 0, 132, 0, 215, 0, 64, 0, 193, 0, 246, 0, 235, 0, 232, 0, 90, 0, 29, 0, 134, 0, 134, 0, 9, 0, 56, 0, 83, 0, 149, 0, 39, 0, 160, 0, 243, 0, 58, 0, 1, 0, 3, 0, 14, 0, 101, 0, 236, 0, 89, 0, 63, 0, 59, 0, 27, 0, 224, 0, 188, 0, 153, 0, 133, 0, 224, 0, 203, 0, 215, 0, 72, 0, 92, 0, 234, 0, 63, 0, 131, 0, 143, 0, 93, 0, 151, 0, 106, 0, 40, 0, 136, 0, 194, 0, 233, 0, 149, 0, 55, 0, 171, 0, 23, 0, 197, 0, 70, 0, 249, 0, 243, 0, 181, 0, 100, 0, 186, 0, 93, 0, 247, 0, 121, 0, 79, 0, 167, 0, 236, 0, 4, 0, 21, 0, 119, 0, 120, 0, 79, 0, 211, 0, 6, 0, 205, 0, 242, 0, 98, 0, 0, 0, 115, 0, 126, 0, 40, 0, 63, 0, 24, 0, 91, 0, 232, 0, 118, 0, 211, 0, 245, 0, 178, 0, 119, 0, 251, 0, 14, 0, 127, 0, 219, 0, 133, 0, 197, 0, 18, 0, 200, 0, 147, 0, 137, 0, 194, 0, 251, 0, 227, 0, 187, 0, 157, 0, 246, 0, 253, 0, 17, 0, 19, 0, 81, 0, 194, 0, 57, 0, 67, 0, 95, 0, 140, 0, 144, 0, 155, 0, 27, 0, 229, 0, 148, 0, 63, 0, 172, 0, 199, 0, 227, 0, 169, 0, 225, 0, 232, 0, 59, 0, 76, 0, 50, 0, 68, 0, 18, 0, 82, 0, 225, 0, 165, 0, 163, 0, 132, 0, 78, 0, 20, 0, 93, 0, 207, 0, 34, 0, 156, 0, 150, 0, 253, 0, 64, 0, 127, 0, 89, 0, 92, 0, 220, 0, 61, 0, 59, 0, 68, 0, 207, 0, 177, 0, 44, 0, 77, 0, 213, 0, 69, 0, 25, 0, 245, 0, 28, 0, 156, 0, 129, 0, 84, 0, 72, 0, 140, 0, 84, 0, 156, 0, 32, 0, 138, 0, 46, 0, 199, 0, 232, 0, 70, 0, 77, 0, 255, 0, 154, 0, 12, 0, 145, 0, 216, 0, 210, 0, 50, 0, 123, 0, 120, 0, 195, 0, 126, 0, 81, 0, 116, 0, 207, 0, 71, 0, 186, 0, 236, 0, 78, 0, 254, 0, 19, 0, 103, 0, 187, 0, 225, 0, 69, 0, 93, 0, 123, 0, 12, 0, 63, 0, 5, 0, 214, 0, 29, 0, 183, 0, 165, 0, 177, 0, 204, 0, 41, 0, 169, 0, 141, 0, 124, 0, 12, 0, 47, 0, 209, 0, 73, 0, 247, 0, 40, 0, 44, 0, 93, 0, 192, 0, 157, 0, 230, 0, 242, 0, 169, 0, 68, 0, 84, 0, 136, 0, 133, 0, 71, 0, 204, 0, 91, 0, 165, 0, 127, 0, 141, 0, 252, 0, 247, 0, 155, 0, 243, 0, 159, 0, 127, 0, 203, 0, 91, 0, 56, 0, 185, 0, 164, 0, 62, 0, 121, 0, 133, 0, 205, 0, 161, 0, 214, 0, 237, 0, 92, 0, 200, 0, 158, 0, 167, 0, 160, 0, 236, 0, 62, 0, 18, 0, 236, 0, 18, 0, 130, 0, 142, 0, 10, 0, 46, 0, 133, 0, 98, 0, 95, 0, 4, 0, 249, 0, 158, 0, 153, 0, 140, 0, 72, 0, 64, 0, 155, 0, 190, 0, 40, 0, 101, 0, 246, 0, 175, 0, 116, 0, 144, 0, 152, 0, 60, 0, 42, 0, 109, 0, 211, 0, 3, 0, 239, 0, 254, 0, 188, 0, 56, 0, 179, 0, 131, 0, 121, 0, 24, 0, 26, 0, 234, 0, 207, 0, 210, 0, 12, 0, 209, 0, 216, 0, 70, 0, 249, 0, 96, 0, 159, 0, 179, 0, 181, 0, 94, 0, 33, 0, 58, 0, 229, 0, 109, 0, 186, 0, 66, 0, 208, 0, 35, 0, 239, 0, 230, 0, 211, 0, 83, 0, 135, 0, 68, 0, 182, 0, 244, 0, 171, 0, 79, 0, 80, 0, 116, 0, 51, 0, 3, 0, 250, 0, 158, 0, 210, 0, 124, 0, 143, 0, 72, 0, 81, 0, 226, 0, 79, 0, 9, 0, 111, 0, 251, 0, 211, 0, 131, 0, 188, 0, 115, 0, 59, 0, 56, 0, 34, 0, 43, 0, 33, 0, 127, 0, 138, 0, 240, 0, 130, 0, 44, 0, 104, 0, 120, 0, 81, 0, 208, 0, 221, 0, 112, 0, 31, 0, 85, 0, 191, 0, 40, 0, 172, 0, 225, 0, 189, 0, 186, 0, 63, 0, 41, 0, 10, 0, 86, 0, 177, 0, 68, 0, 199, 0, 27, 0, 221, 0, 49, 0, 130, 0, 155, 0, 40, 0, 123, 0, 55, 0, 156, 0, 88, 0, 201, 0, 186, 0, 218, 0, 110, 0, 233, 0, 24, 0, 39, 0, 208, 0, 246, 0, 59, 0, 110, 0, 83, 0, 132, 0, 87, 0, 23, 0, 182, 0, 214, 0, 39, 0, 135, 0, 43, 0, 139, 0, 11, 0, 86, 0, 97, 0, 151, 0, 67, 0, 17, 0, 113, 0, 214, 0, 47, 0, 198, 0, 191, 0, 119, 0, 69, 0, 32, 0, 0, 0, 194, 0, 127, 0, 189, 0, 85, 0, 238, 0, 166, 0, 205, 0, 125, 0, 79, 0, 88, 0, 56, 0, 166, 0, 240, 0, 28, 0, 253, 0, 40, 0, 251, 0, 5, 0, 232, 0, 237, 0, 86, 0, 144, 0, 16, 0, 190, 0, 33, 0, 152, 0, 246, 0, 249, 0, 40, 0, 166, 0, 72, 0, 35, 0, 192, 0, 147, 0, 229, 0, 218, 0, 137, 0, 37, 0, 130, 0, 136, 0, 187, 0, 14, 0, 211, 0, 193, 0, 184, 0, 168, 0, 213, 0, 8, 0, 30, 0, 0, 0, 6, 0, 136, 0, 54, 0, 174, 0, 148, 0, 86, 0, 154, 0, 177, 0, 24, 0, 2, 0, 234, 0, 48, 0, 3, 0, 78, 0, 84, 0, 22, 0, 123, 0, 40, 0, 171, 0, 228, 0, 19, 0, 1, 0, 14, 0, 113, 0, 229, 0, 69, 0, 23, 0, 141, 0, 20, 0, 160, 0, 67, 0, 50, 0, 157, 0, 49, 0, 69, 0, 57, 0, 126, 0, 238, 0, 12, 0, 185, 0, 254, 0, 162, 0, 26, 0, 89, 0, 223, 0, 49, 0, 233, 0, 15, 0, 135, 0, 89, 0, 30, 0, 99, 0, 101, 0, 184, 0, 141, 0, 194, 0, 98, 0, 147, 0, 238, 0, 117, 0, 13, 0, 156, 0, 24, 0, 138, 0, 199, 0, 121, 0, 186, 0, 15, 0, 234, 0, 111, 0, 84, 0, 96, 0, 45, 0, 195, 0, 171, 0, 41, 0, 153, 0, 54, 0, 173, 0, 235, 0, 204, 0, 221, 0, 88, 0, 233, 0, 65, 0, 208, 0, 120, 0, 206, 0, 252, 0, 82, 0, 185, 0, 44, 0, 48, 0, 198, 0, 155, 0, 17, 0, 155, 0, 121, 0, 70, 0, 13, 0, 148, 0, 23, 0, 148, 0, 94, 0, 232, 0, 72, 0, 27, 0, 166, 0, 185, 0, 200, 0, 118, 0, 115, 0, 200, 0, 182, 0);
    signal scenario_full  : scenario_type := (176, 31, 66, 31, 159, 31, 63, 31, 164, 31, 33, 31, 114, 31, 93, 31, 199, 31, 84, 31, 160, 31, 237, 31, 44, 31, 21, 31, 80, 31, 80, 30, 115, 31, 113, 31, 229, 31, 132, 31, 171, 31, 6, 31, 202, 31, 44, 31, 173, 31, 144, 31, 212, 31, 51, 31, 15, 31, 173, 31, 140, 31, 126, 31, 12, 31, 252, 31, 195, 31, 254, 31, 249, 31, 215, 31, 17, 31, 180, 31, 33, 31, 163, 31, 186, 31, 207, 31, 16, 31, 200, 31, 157, 31, 48, 31, 214, 31, 87, 31, 118, 31, 71, 31, 18, 31, 13, 31, 13, 31, 177, 31, 80, 31, 56, 31, 20, 31, 73, 31, 24, 31, 29, 31, 214, 31, 82, 31, 191, 31, 191, 30, 195, 31, 254, 31, 40, 31, 222, 31, 170, 31, 123, 31, 215, 31, 189, 31, 146, 31, 132, 31, 71, 31, 208, 31, 203, 31, 193, 31, 234, 31, 1, 31, 245, 31, 117, 31, 23, 31, 23, 30, 113, 31, 121, 31, 26, 31, 79, 31, 223, 31, 137, 31, 209, 31, 64, 31, 252, 31, 9, 31, 13, 31, 226, 31, 2, 31, 42, 31, 174, 31, 122, 31, 219, 31, 219, 31, 33, 31, 239, 31, 179, 31, 122, 31, 64, 31, 13, 31, 72, 31, 125, 31, 205, 31, 162, 31, 59, 31, 113, 31, 43, 31, 63, 31, 224, 31, 14, 31, 94, 31, 33, 31, 66, 31, 20, 31, 49, 31, 160, 31, 52, 31, 34, 31, 9, 31, 253, 31, 27, 31, 14, 31, 135, 31, 109, 31, 204, 31, 121, 31, 237, 31, 171, 31, 173, 31, 112, 31, 133, 31, 247, 31, 81, 31, 35, 31, 73, 31, 129, 31, 152, 31, 193, 31, 92, 31, 74, 31, 45, 31, 12, 31, 54, 31, 36, 31, 224, 31, 93, 31, 84, 31, 37, 31, 39, 31, 188, 31, 245, 31, 112, 31, 239, 31, 243, 31, 14, 31, 135, 31, 225, 31, 78, 31, 103, 31, 34, 31, 34, 30, 6, 31, 81, 31, 254, 31, 11, 31, 121, 31, 217, 31, 119, 31, 39, 31, 130, 31, 190, 31, 18, 31, 145, 31, 190, 31, 72, 31, 251, 31, 222, 31, 172, 31, 200, 31, 136, 31, 120, 31, 37, 31, 86, 31, 125, 31, 160, 31, 94, 31, 222, 31, 146, 31, 146, 31, 221, 31, 66, 31, 247, 31, 129, 31, 150, 31, 188, 31, 67, 31, 19, 31, 128, 31, 158, 31, 146, 31, 206, 31, 99, 31, 48, 31, 220, 31, 3, 31, 173, 31, 67, 31, 3, 31, 126, 31, 203, 31, 234, 31, 81, 31, 81, 30, 11, 31, 227, 31, 162, 31, 38, 31, 156, 31, 17, 31, 95, 31, 202, 31, 209, 31, 145, 31, 134, 31, 57, 31, 136, 31, 159, 31, 103, 31, 37, 31, 12, 31, 209, 31, 187, 31, 219, 31, 177, 31, 244, 31, 121, 31, 220, 31, 59, 31, 91, 31, 155, 31, 119, 31, 58, 31, 115, 31, 235, 31, 67, 31, 79, 31, 28, 31, 107, 31, 7, 31, 120, 31, 7, 31, 131, 31, 204, 31, 77, 31, 158, 31, 201, 31, 120, 31, 168, 31, 110, 31, 81, 31, 238, 31, 189, 31, 188, 31, 67, 31, 51, 31, 185, 31, 153, 31, 219, 31, 35, 31, 192, 31, 149, 31, 110, 31, 97, 31, 227, 31, 67, 31, 245, 31, 138, 31, 99, 31, 7, 31, 189, 31, 51, 31, 185, 31, 185, 30, 235, 31, 56, 31, 245, 31, 46, 31, 233, 31, 54, 31, 179, 31, 95, 31, 221, 31, 78, 31, 253, 31, 183, 31, 229, 31, 119, 31, 67, 31, 172, 31, 58, 31, 16, 31, 166, 31, 150, 31, 192, 31, 54, 31, 234, 31, 176, 31, 96, 31, 175, 31, 106, 31, 181, 31, 48, 31, 85, 31, 202, 31, 154, 31, 151, 31, 66, 31, 104, 31, 28, 31, 244, 31, 76, 31, 183, 31, 254, 31, 150, 31, 117, 31, 243, 31, 153, 31, 65, 31, 184, 31, 30, 31, 177, 31, 245, 31, 225, 31, 255, 31, 173, 31, 127, 31, 163, 31, 204, 31, 59, 31, 68, 31, 76, 31, 181, 31, 96, 31, 131, 31, 14, 31, 242, 31, 35, 31, 31, 31, 195, 31, 145, 31, 153, 31, 12, 31, 180, 31, 175, 31, 248, 31, 73, 31, 100, 31, 4, 31, 186, 31, 14, 31, 170, 31, 194, 31, 102, 31, 118, 31, 252, 31, 191, 31, 175, 31, 245, 31, 182, 31, 75, 31, 210, 31, 41, 31, 177, 31, 101, 31, 149, 31, 9, 31, 119, 31, 30, 31, 49, 31, 119, 31, 164, 31, 118, 31, 245, 31, 105, 31, 92, 31, 201, 31, 175, 31, 167, 31, 224, 31, 99, 31, 14, 31, 63, 31, 104, 31, 189, 31, 174, 31, 84, 31, 160, 31, 206, 31, 4, 31, 20, 31, 173, 31, 187, 31, 82, 31, 46, 31, 234, 31, 217, 31, 20, 31, 47, 31, 8, 31, 119, 31, 31, 31, 198, 31, 25, 31, 170, 31, 139, 31, 218, 31, 4, 31, 207, 31, 65, 31, 222, 31, 132, 31, 215, 31, 64, 31, 193, 31, 246, 31, 235, 31, 232, 31, 90, 31, 29, 31, 134, 31, 134, 31, 9, 31, 56, 31, 83, 31, 149, 31, 39, 31, 160, 31, 243, 31, 58, 31, 1, 31, 3, 31, 14, 31, 101, 31, 236, 31, 89, 31, 63, 31, 59, 31, 27, 31, 224, 31, 188, 31, 153, 31, 133, 31, 224, 31, 203, 31, 215, 31, 72, 31, 92, 31, 234, 31, 63, 31, 131, 31, 143, 31, 93, 31, 151, 31, 106, 31, 40, 31, 136, 31, 194, 31, 233, 31, 149, 31, 55, 31, 171, 31, 23, 31, 197, 31, 70, 31, 249, 31, 243, 31, 181, 31, 100, 31, 186, 31, 93, 31, 247, 31, 121, 31, 79, 31, 167, 31, 236, 31, 4, 31, 21, 31, 119, 31, 120, 31, 79, 31, 211, 31, 6, 31, 205, 31, 242, 31, 98, 31, 98, 30, 115, 31, 126, 31, 40, 31, 63, 31, 24, 31, 91, 31, 232, 31, 118, 31, 211, 31, 245, 31, 178, 31, 119, 31, 251, 31, 14, 31, 127, 31, 219, 31, 133, 31, 197, 31, 18, 31, 200, 31, 147, 31, 137, 31, 194, 31, 251, 31, 227, 31, 187, 31, 157, 31, 246, 31, 253, 31, 17, 31, 19, 31, 81, 31, 194, 31, 57, 31, 67, 31, 95, 31, 140, 31, 144, 31, 155, 31, 27, 31, 229, 31, 148, 31, 63, 31, 172, 31, 199, 31, 227, 31, 169, 31, 225, 31, 232, 31, 59, 31, 76, 31, 50, 31, 68, 31, 18, 31, 82, 31, 225, 31, 165, 31, 163, 31, 132, 31, 78, 31, 20, 31, 93, 31, 207, 31, 34, 31, 156, 31, 150, 31, 253, 31, 64, 31, 127, 31, 89, 31, 92, 31, 220, 31, 61, 31, 59, 31, 68, 31, 207, 31, 177, 31, 44, 31, 77, 31, 213, 31, 69, 31, 25, 31, 245, 31, 28, 31, 156, 31, 129, 31, 84, 31, 72, 31, 140, 31, 84, 31, 156, 31, 32, 31, 138, 31, 46, 31, 199, 31, 232, 31, 70, 31, 77, 31, 255, 31, 154, 31, 12, 31, 145, 31, 216, 31, 210, 31, 50, 31, 123, 31, 120, 31, 195, 31, 126, 31, 81, 31, 116, 31, 207, 31, 71, 31, 186, 31, 236, 31, 78, 31, 254, 31, 19, 31, 103, 31, 187, 31, 225, 31, 69, 31, 93, 31, 123, 31, 12, 31, 63, 31, 5, 31, 214, 31, 29, 31, 183, 31, 165, 31, 177, 31, 204, 31, 41, 31, 169, 31, 141, 31, 124, 31, 12, 31, 47, 31, 209, 31, 73, 31, 247, 31, 40, 31, 44, 31, 93, 31, 192, 31, 157, 31, 230, 31, 242, 31, 169, 31, 68, 31, 84, 31, 136, 31, 133, 31, 71, 31, 204, 31, 91, 31, 165, 31, 127, 31, 141, 31, 252, 31, 247, 31, 155, 31, 243, 31, 159, 31, 127, 31, 203, 31, 91, 31, 56, 31, 185, 31, 164, 31, 62, 31, 121, 31, 133, 31, 205, 31, 161, 31, 214, 31, 237, 31, 92, 31, 200, 31, 158, 31, 167, 31, 160, 31, 236, 31, 62, 31, 18, 31, 236, 31, 18, 31, 130, 31, 142, 31, 10, 31, 46, 31, 133, 31, 98, 31, 95, 31, 4, 31, 249, 31, 158, 31, 153, 31, 140, 31, 72, 31, 64, 31, 155, 31, 190, 31, 40, 31, 101, 31, 246, 31, 175, 31, 116, 31, 144, 31, 152, 31, 60, 31, 42, 31, 109, 31, 211, 31, 3, 31, 239, 31, 254, 31, 188, 31, 56, 31, 179, 31, 131, 31, 121, 31, 24, 31, 26, 31, 234, 31, 207, 31, 210, 31, 12, 31, 209, 31, 216, 31, 70, 31, 249, 31, 96, 31, 159, 31, 179, 31, 181, 31, 94, 31, 33, 31, 58, 31, 229, 31, 109, 31, 186, 31, 66, 31, 208, 31, 35, 31, 239, 31, 230, 31, 211, 31, 83, 31, 135, 31, 68, 31, 182, 31, 244, 31, 171, 31, 79, 31, 80, 31, 116, 31, 51, 31, 3, 31, 250, 31, 158, 31, 210, 31, 124, 31, 143, 31, 72, 31, 81, 31, 226, 31, 79, 31, 9, 31, 111, 31, 251, 31, 211, 31, 131, 31, 188, 31, 115, 31, 59, 31, 56, 31, 34, 31, 43, 31, 33, 31, 127, 31, 138, 31, 240, 31, 130, 31, 44, 31, 104, 31, 120, 31, 81, 31, 208, 31, 221, 31, 112, 31, 31, 31, 85, 31, 191, 31, 40, 31, 172, 31, 225, 31, 189, 31, 186, 31, 63, 31, 41, 31, 10, 31, 86, 31, 177, 31, 68, 31, 199, 31, 27, 31, 221, 31, 49, 31, 130, 31, 155, 31, 40, 31, 123, 31, 55, 31, 156, 31, 88, 31, 201, 31, 186, 31, 218, 31, 110, 31, 233, 31, 24, 31, 39, 31, 208, 31, 246, 31, 59, 31, 110, 31, 83, 31, 132, 31, 87, 31, 23, 31, 182, 31, 214, 31, 39, 31, 135, 31, 43, 31, 139, 31, 11, 31, 86, 31, 97, 31, 151, 31, 67, 31, 17, 31, 113, 31, 214, 31, 47, 31, 198, 31, 191, 31, 119, 31, 69, 31, 32, 31, 32, 30, 194, 31, 127, 31, 189, 31, 85, 31, 238, 31, 166, 31, 205, 31, 125, 31, 79, 31, 88, 31, 56, 31, 166, 31, 240, 31, 28, 31, 253, 31, 40, 31, 251, 31, 5, 31, 232, 31, 237, 31, 86, 31, 144, 31, 16, 31, 190, 31, 33, 31, 152, 31, 246, 31, 249, 31, 40, 31, 166, 31, 72, 31, 35, 31, 192, 31, 147, 31, 229, 31, 218, 31, 137, 31, 37, 31, 130, 31, 136, 31, 187, 31, 14, 31, 211, 31, 193, 31, 184, 31, 168, 31, 213, 31, 8, 31, 30, 31, 30, 30, 6, 31, 136, 31, 54, 31, 174, 31, 148, 31, 86, 31, 154, 31, 177, 31, 24, 31, 2, 31, 234, 31, 48, 31, 3, 31, 78, 31, 84, 31, 22, 31, 123, 31, 40, 31, 171, 31, 228, 31, 19, 31, 1, 31, 14, 31, 113, 31, 229, 31, 69, 31, 23, 31, 141, 31, 20, 31, 160, 31, 67, 31, 50, 31, 157, 31, 49, 31, 69, 31, 57, 31, 126, 31, 238, 31, 12, 31, 185, 31, 254, 31, 162, 31, 26, 31, 89, 31, 223, 31, 49, 31, 233, 31, 15, 31, 135, 31, 89, 31, 30, 31, 99, 31, 101, 31, 184, 31, 141, 31, 194, 31, 98, 31, 147, 31, 238, 31, 117, 31, 13, 31, 156, 31, 24, 31, 138, 31, 199, 31, 121, 31, 186, 31, 15, 31, 234, 31, 111, 31, 84, 31, 96, 31, 45, 31, 195, 31, 171, 31, 41, 31, 153, 31, 54, 31, 173, 31, 235, 31, 204, 31, 221, 31, 88, 31, 233, 31, 65, 31, 208, 31, 120, 31, 206, 31, 252, 31, 82, 31, 185, 31, 44, 31, 48, 31, 198, 31, 155, 31, 17, 31, 155, 31, 121, 31, 70, 31, 13, 31, 148, 31, 23, 31, 148, 31, 94, 31, 232, 31, 72, 31, 27, 31, 166, 31, 185, 31, 200, 31, 118, 31, 115, 31, 200, 31, 182, 31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
